library verilog;
use verilog.vl_types.all;
entity FFT_vlg_vec_tst is
end FFT_vlg_vec_tst;
