-----------------------------------------------------------
--
-- Copyright (c) 2020, nmrenyi <ry18@mails.tsinghua.edu.cn>
-- Referenced to https://github.com/Ugon/fpga-fft-equalizer
-----------------------------------------------------------
-- fft_utils.vhd
-- create time: 2020-05-01
-- target chip: EP2C70F672C8
-- main function: functions used in the project.
-----------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.fft_twiddle_factors_64.all;

package fft_utils is
	constant tw_size: integer := tw_size;

	procedure complex_twiddle_mult(
		twiddle_num:  in  integer;
		fft_size_exp: in  integer;
		in_re:  	  in  signed;
		in_im:  	  in  signed;
		out_re: 	  out signed;
		out_im: 	  out signed);

	function bit_reverse(number: unsigned) return unsigned;

	function bit_reverse(number: std_logic_vector) return std_logic_vector;

	function negate_all(samples: std_logic_vector; number_of_samples: integer; bits_per_sample: integer) return std_logic_vector;

	function shuffle(samples: std_logic_vector; fft_size_exp: integer; bits_per_sample: integer) return std_logic_vector;
	
	function divide_and_resize_all(samples: std_logic_vector; number_of_samples: integer; old_bits_per_sample: integer; divisor: integer; new_bits_per_sample: integer) return std_logic_vector;

	function resize_all(samples: std_logic_vector; number_of_samples: integer; old_bits_per_sample: integer; new_bits_per_sample: integer) return std_logic_vector;

end;

package body fft_utils is

	procedure complex_twiddle_mult(
		twiddle_num:  in  integer;
		fft_size_exp: in  integer;
		in_re:        in  signed;
		in_im:        in  signed;
		out_re:       out signed;
		out_im:       out signed)
	is
		constant tw_re:         signed(tw_size - 1 downto 0) := re_64(twiddle_num * 2**(tw_array_size_exp - fft_size_exp));
		constant tw_im:         signed(tw_size - 1 downto 0) := im_64(twiddle_num * 2**(tw_array_size_exp - fft_size_exp));

		variable multed1:       signed(in_re'length + tw_re'length - 1 downto 0);
		variable multed2:       signed(in_im'length + tw_im'length - 1 downto 0);
		variable multed3:       signed(in_re'length + tw_im'length - 1 downto 0);
		variable multed4:       signed(in_im'length + tw_re'length - 1 downto 0);

		variable multed1_trunc: signed(in_re'length - 1 downto 0);
		variable multed2_trunc: signed(in_im'length - 1 downto 0);
		variable multed3_trunc: signed(in_re'length - 1 downto 0);
		variable multed4_trunc: signed(in_im'length - 1 downto 0);

	begin
		if twiddle_num = 0 then
			out_re := in_re;  
			out_im := in_im;  
		elsif twiddle_num * 2**(8 - fft_size_exp) = 64 then
			out_re := - in_im;  
			out_im :=   in_re;
		else
			multed1 := in_re * tw_re;
			multed2 := in_im * tw_im;
			multed3 := in_re * tw_im;
			multed4 := in_im * tw_re;

			multed1_trunc := multed1(multed1'length - 2 downto tw_size - 1);
			multed2_trunc := multed2(multed2'length - 2 downto tw_size - 1);
			multed3_trunc := multed3(multed3'length - 2 downto tw_size - 1);
			multed4_trunc := multed4(multed4'length - 2 downto tw_size - 1);

			out_re := multed1_trunc - multed2_trunc;
			out_im := multed3_trunc + multed4_trunc;
		end if;

	end complex_twiddle_mult;

	function bit_reverse(number: unsigned) return unsigned is
		variable reversed: unsigned(number'range);
		alias number_alias: unsigned(number'reverse_range) is number;
	begin
		for i in number_alias'range loop
			reversed(i) := number_alias(i);
		end loop;
		return reversed;
	end function;

	function bit_reverse(number: std_logic_vector) return std_logic_vector is
		variable reversed: std_logic_vector(number'range);
		alias number_alias: std_logic_vector(number'reverse_range) is number;
	begin
		for i in number_alias'range loop
			reversed(i) := number_alias(i);
		end loop;
		return reversed;
	end function;

	function negate_all(samples: std_logic_vector; number_of_samples: integer; bits_per_sample: integer) return std_logic_vector is
		variable negated: std_logic_vector(samples'length - 1 downto 0);
	begin
		for i in number_of_samples - 1 downto 0 loop
			negated((i + 1) * bits_per_sample - 1 downto i * bits_per_sample) := std_logic_vector(- signed(samples((i + 1) * bits_per_sample - 1 downto i * bits_per_sample)));
		end loop;
		return negated;
	end function;

	function shuffle(samples: std_logic_vector; fft_size_exp: integer; bits_per_sample: integer) return std_logic_vector is
		variable shuffled:  std_logic_vector(samples'length - 1 downto 0);
		variable reversed_i: integer;
	begin
		for i in 2**fft_size_exp - 1 downto 0 loop
			reversed_i := to_integer(bit_reverse(to_unsigned(i, fft_size_exp)));
			shuffled((reversed_i + 1) * bits_per_sample - 1 downto reversed_i * bits_per_sample) := std_logic_vector(signed(samples((i + 1) * bits_per_sample - 1 downto i * bits_per_sample)));
		end loop;
		return shuffled;
	end function;

	function divide_and_resize_all(samples: std_logic_vector; number_of_samples: integer; old_bits_per_sample: integer; divisor: integer; new_bits_per_sample: integer) return std_logic_vector is
		variable output_vector: std_logic_vector(number_of_samples * new_bits_per_sample - 1 downto 0);
	begin
		for i in number_of_samples - 1 downto 0 loop
			output_vector((i + 1) * (new_bits_per_sample) - 1 downto i * (new_bits_per_sample))
				:= std_logic_vector(resize(signed(samples((i + 1) * old_bits_per_sample - 1 downto i * old_bits_per_sample)) / divisor, new_bits_per_sample));
		end loop;
		return output_vector;
	end function;

	function resize_all(samples: std_logic_vector; number_of_samples: integer; old_bits_per_sample: integer; new_bits_per_sample: integer) return std_logic_vector is
		variable output_vector: std_logic_vector(number_of_samples * new_bits_per_sample - 1 downto 0);
	begin
		for i in number_of_samples - 1 downto 0 loop
			output_vector((i + 1) * (new_bits_per_sample) - 1 downto i * (new_bits_per_sample))
				:= std_logic_vector(resize(signed(samples((i + 1) * old_bits_per_sample - 1 downto i * old_bits_per_sample)), new_bits_per_sample));
		end loop;
		return output_vector;
	end function;

end package body;