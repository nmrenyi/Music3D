-- library ieee;
-- use ieee.std_logic_1164.all;
-- use ieee.numeric_std.all;

-- package fft_twiddle_factors_64 is
-- 	constant tw_size:           integer := 16;
-- 	constant tw_array_size_exp: integer := 6;
	
-- 	type arr is array (0 to 2**(tw_array_size_exp - 1) - 1) of signed(tw_size - 1 downto 0);

-- 	constant re_64: arr := (
-- 		0 =>  "0111111111111111", --'one' 16-bit approximation
-- 		1 =>  "0111111101100010",
-- 		2 =>  "0111110110001010",
-- 		3 =>  "0111101001111101",
-- 		4 =>  "0111011001000010",
-- 		5 =>  "0111000011100011",
-- 		6 =>  "0110101001101110",
-- 		7 =>  "0110001011110010",
-- 		8 =>  "0101101010000010",
-- 		9 =>  "0101000100110100",
-- 		10 => "0100011100011101",
-- 		11 => "0011110001010111",
-- 		12 => "0011000011111100",
-- 		13 => "0010010100101000",
-- 		14 => "0001100011111001",
-- 		15 => "0000110010001100",
-- 		16 => "0000000000000000",
-- 		17 => "1111001101110100",
-- 		18 => "1110011100000111",
-- 		19 => "1101101011011000",
-- 		20 => "1100111100000100",
-- 		21 => "1100001110101001",
-- 		22 => "1011100011100011",
-- 		23 => "1010111011001100",
-- 		24 => "1010010101111110",
-- 		25 => "1001110100001110",
-- 		26 => "1001010110010010",
-- 		27 => "1000111100011101",
-- 		28 => "1000100110111110",
-- 		29 => "1000010110000011",
-- 		30 => "1000001001110110",
-- 		31 => "1000000010011110");

-- 	constant im_64: arr := (
-- 		0 =>  "0000000000000000",
-- 		1 =>  "0000110010001100",
-- 		2 =>  "0001100011111001",
-- 		3 =>  "0010010100101000",
-- 		4 =>  "0011000011111100",
-- 		5 =>  "0011110001010111",
-- 		6 =>  "0100011100011101",
-- 		7 =>  "0101000100110100",
-- 		8 =>  "0101101010000010",
-- 		9 =>  "0110001011110010",
-- 		10 => "0110101001101110",
-- 		11 => "0111000011100011",
-- 		12 => "0111011001000010",
-- 		13 => "0111101001111101",
-- 		14 => "0111110110001010",
-- 		15 => "0111111101100010",
-- 		16 => "0111111111111111", --'one' 16-bit approximation
-- 		17 => "0111111101100010",
-- 		18 => "0111110110001010",
-- 		19 => "0111101001111101",
-- 		20 => "0111011001000010",
-- 		21 => "0111000011100011",
-- 		22 => "0110101001101110",
-- 		23 => "0110001011110010",
-- 		24 => "0101101010000010",
-- 		25 => "0101000100110100",
-- 		26 => "0100011100011101",
-- 		27 => "0011110001010111",
-- 		28 => "0011000011111100",
-- 		29 => "0010010100101000",
-- 		30 => "0001100011111001",
-- 		31 => "0000110010001100");
-- end;




library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fft_twiddle_factors_64 is
	constant tw_size:           integer := 16;
	constant tw_array_size_exp: integer := 10;
	
	type arr is array (0 to 2**(tw_array_size_exp - 1) - 1) of signed(tw_size - 1 downto 0);

	constant re_64: arr := (
		0 => "0111111111111111",
		1 => "0111111111111110",
		2 => "0111111111111100",
		3 => "0111111111111001",
		4 => "0111111111110101",
		5 => "0111111111101111",
		6 => "0111111111101000",
		7 => "0111111111100000",
		8 => "0111111111010111",
		9 => "0111111111001101",
		10 => "0111111111000001",
		11 => "0111111110110100",
		12 => "0111111110100110",
		13 => "0111111110010110",
		14 => "0111111110000110",
		15 => "0111111101110100",
		16 => "0111111101100001",
		17 => "0111111101001100",
		18 => "0111111100110111",
		19 => "0111111100100000",
		20 => "0111111100001000",
		21 => "0111111011101111",
		22 => "0111111011010100",
		23 => "0111111010111001",
		24 => "0111111010011100",
		25 => "0111111001111110",
		26 => "0111111001011110",
		27 => "0111111000111110",
		28 => "0111111000011100",
		29 => "0111110111111001",
		30 => "0111110111010101",
		31 => "0111110110110000",
		32 => "0111110110001001",
		33 => "0111110101100001",
		34 => "0111110100111000",
		35 => "0111110100001110",
		36 => "0111110011100010",
		37 => "0111110010110110",
		38 => "0111110010001000",
		39 => "0111110001011001",
		40 => "0111110000101001",
		41 => "0111101111110111",
		42 => "0111101111000100",
		43 => "0111101110010001",
		44 => "0111101101011100",
		45 => "0111101100100101",
		46 => "0111101011101110",
		47 => "0111101010110101",
		48 => "0111101001111100",
		49 => "0111101001000001",
		50 => "0111101000000100",
		51 => "0111100111000111",
		52 => "0111100110001001",
		53 => "0111100101001001",
		54 => "0111100100001000",
		55 => "0111100011000110",
		56 => "0111100010000011",
		57 => "0111100000111111",
		58 => "0111011111111001",
		59 => "0111011110110011",
		60 => "0111011101101011",
		61 => "0111011100100010",
		62 => "0111011011011000",
		63 => "0111011010001101",
		64 => "0111011001000000",
		65 => "0111010111110011",
		66 => "0111010110100100",
		67 => "0111010101010100",
		68 => "0111010100000011",
		69 => "0111010010110001",
		70 => "0111010001011110",
		71 => "0111010000001010",
		72 => "0111001110110101",
		73 => "0111001101011110",
		74 => "0111001100000110",
		75 => "0111001010101110",
		76 => "0111001001010100",
		77 => "0111000111111001",
		78 => "0111000110011101",
		79 => "0111000101000000",
		80 => "0111000011100001",
		81 => "0111000010000010",
		82 => "0111000000100010",
		83 => "0110111111000000",
		84 => "0110111101011110",
		85 => "0110111011111010",
		86 => "0110111010010101",
		87 => "0110111000110000",
		88 => "0110110111001001",
		89 => "0110110101100001",
		90 => "0110110011111000",
		91 => "0110110010001110",
		92 => "0110110000100011",
		93 => "0110101110110111",
		94 => "0110101101001010",
		95 => "0110101011011011",
		96 => "0110101001101100",
		97 => "0110100111111100",
		98 => "0110100110001011",
		99 => "0110100100011001",
		100 => "0110100010100101",
		101 => "0110100000110001",
		102 => "0110011110111100",
		103 => "0110011101000101",
		104 => "0110011011001110",
		105 => "0110011001010110",
		106 => "0110010111011101",
		107 => "0110010101100010",
		108 => "0110010011100111",
		109 => "0110010001101011",
		110 => "0110001111101110",
		111 => "0110001101110000",
		112 => "0110001011110001",
		113 => "0110001001110001",
		114 => "0110000111110000",
		115 => "0110000101101110",
		116 => "0110000011101011",
		117 => "0110000001100111",
		118 => "0101111111100010",
		119 => "0101111101011101",
		120 => "0101111011010110",
		121 => "0101111001001111",
		122 => "0101110111000110",
		123 => "0101110100111101",
		124 => "0101110010110011",
		125 => "0101110000101000",
		126 => "0101101110011100",
		127 => "0101101100001111",
		128 => "0101101010000001",
		129 => "0101100111110011",
		130 => "0101100101100011",
		131 => "0101100011010011",
		132 => "0101100001000010",
		133 => "0101011110110000",
		134 => "0101011100011101",
		135 => "0101011010001001",
		136 => "0101010111110100",
		137 => "0101010101011111",
		138 => "0101010011001001",
		139 => "0101010000110010",
		140 => "0101001110011010",
		141 => "0101001100000001",
		142 => "0101001001101000",
		143 => "0101000111001110",
		144 => "0101000100110011",
		145 => "0101000010010111",
		146 => "0100111111111010",
		147 => "0100111101011101",
		148 => "0100111010111111",
		149 => "0100111000100000",
		150 => "0100110110000000",
		151 => "0100110011100000",
		152 => "0100110000111111",
		153 => "0100101110011101",
		154 => "0100101011111010",
		155 => "0100101001010111",
		156 => "0100100110110011",
		157 => "0100100100001110",
		158 => "0100100001101001",
		159 => "0100011111000011",
		160 => "0100011100011100",
		161 => "0100011001110100",
		162 => "0100010111001100",
		163 => "0100010100100011",
		164 => "0100010001111010",
		165 => "0100001111010000",
		166 => "0100001100100101",
		167 => "0100001001111001",
		168 => "0100000111001101",
		169 => "0100000100100000",
		170 => "0100000001110011",
		171 => "0011111111000101",
		172 => "0011111100010110",
		173 => "0011111001100111",
		174 => "0011110110110111",
		175 => "0011110100000111",
		176 => "0011110001010110",
		177 => "0011101110100100",
		178 => "0011101011110010",
		179 => "0011101000111111",
		180 => "0011100110001100",
		181 => "0011100011011000",
		182 => "0011100000100100",
		183 => "0011011101101111",
		184 => "0011011010111001",
		185 => "0011011000000011",
		186 => "0011010101001101",
		187 => "0011010010010110",
		188 => "0011001111011110",
		189 => "0011001100100110",
		190 => "0011001001101101",
		191 => "0011000110110100",
		192 => "0011000011111011",
		193 => "0011000001000001",
		194 => "0010111110000110",
		195 => "0010111011001100",
		196 => "0010111000010000",
		197 => "0010110101010100",
		198 => "0010110010011000",
		199 => "0010101111011011",
		200 => "0010101100011110",
		201 => "0010101001100001",
		202 => "0010100110100011",
		203 => "0010100011100101",
		204 => "0010100000100110",
		205 => "0010011101100111",
		206 => "0010011010100111",
		207 => "0010010111100111",
		208 => "0010010100100111",
		209 => "0010010001100111",
		210 => "0010001110100110",
		211 => "0010001011100100",
		212 => "0010001000100011",
		213 => "0010000101100001",
		214 => "0010000010011111",
		215 => "0001111111011100",
		216 => "0001111100011001",
		217 => "0001111001010110",
		218 => "0001110110010011",
		219 => "0001110011001111",
		220 => "0001110000001011",
		221 => "0001101101000110",
		222 => "0001101010000010",
		223 => "0001100110111101",
		224 => "0001100011111000",
		225 => "0001100000110011",
		226 => "0001011101101101",
		227 => "0001011010100111",
		228 => "0001010111100001",
		229 => "0001010100011011",
		230 => "0001010001010101",
		231 => "0001001110001110",
		232 => "0001001011000111",
		233 => "0001001000000000",
		234 => "0001000100111001",
		235 => "0001000001110010",
		236 => "0000111110101011",
		237 => "0000111011100011",
		238 => "0000111000011011",
		239 => "0000110101010011",
		240 => "0000110010001011",
		241 => "0000101111000011",
		242 => "0000101011111011",
		243 => "0000101000110010",
		244 => "0000100101101010",
		245 => "0000100010100001",
		246 => "0000011111011001",
		247 => "0000011100010000",
		248 => "0000011001000111",
		249 => "0000010101111110",
		250 => "0000010010110110",
		251 => "0000001111101101",
		252 => "0000001100100100",
		253 => "0000001001011011",
		254 => "0000000110010010",
		255 => "0000000011001001",
		256 => "0000000000000000",
		257 => "1111111100110110",
		258 => "1111111001101101",
		259 => "1111110110100100",
		260 => "1111110011011011",
		261 => "1111110000010010",
		262 => "1111101101001001",
		263 => "1111101010000001",
		264 => "1111100110111000",
		265 => "1111100011101111",
		266 => "1111100000100110",
		267 => "1111011101011110",
		268 => "1111011010010101",
		269 => "1111010111001101",
		270 => "1111010100000100",
		271 => "1111010000111100",
		272 => "1111001101110100",
		273 => "1111001010101100",
		274 => "1111000111100100",
		275 => "1111000100011100",
		276 => "1111000001010100",
		277 => "1110111110001101",
		278 => "1110111011000110",
		279 => "1110110111111111",
		280 => "1110110100111000",
		281 => "1110110001110001",
		282 => "1110101110101010",
		283 => "1110101011100100",
		284 => "1110101000011110",
		285 => "1110100101011000",
		286 => "1110100010010010",
		287 => "1110011111001100",
		288 => "1110011100000111",
		289 => "1110011001000010",
		290 => "1110010101111101",
		291 => "1110010010111001",
		292 => "1110001111110100",
		293 => "1110001100110000",
		294 => "1110001001101100",
		295 => "1110000110101001",
		296 => "1110000011100110",
		297 => "1110000000100011",
		298 => "1101111101100000",
		299 => "1101111010011110",
		300 => "1101110111011100",
		301 => "1101110100011011",
		302 => "1101110001011001",
		303 => "1101101110011000",
		304 => "1101101011011000",
		305 => "1101101000011000",
		306 => "1101100101011000",
		307 => "1101100010011000",
		308 => "1101011111011001",
		309 => "1101011100011010",
		310 => "1101011001011100",
		311 => "1101010110011110",
		312 => "1101010011100001",
		313 => "1101010000100100",
		314 => "1101001101100111",
		315 => "1101001010101011",
		316 => "1101000111101111",
		317 => "1101000100110011",
		318 => "1101000001111001",
		319 => "1100111110111110",
		320 => "1100111100000100",
		321 => "1100111001001011",
		322 => "1100110110010010",
		323 => "1100110011011001",
		324 => "1100110000100001",
		325 => "1100101101101001",
		326 => "1100101010110010",
		327 => "1100100111111100",
		328 => "1100100101000110",
		329 => "1100100010010000",
		330 => "1100011111011011",
		331 => "1100011100100111",
		332 => "1100011001110011",
		333 => "1100010111000000",
		334 => "1100010100001101",
		335 => "1100010001011011",
		336 => "1100001110101001",
		337 => "1100001011111000",
		338 => "1100001001001000",
		339 => "1100000110011000",
		340 => "1100000011101001",
		341 => "1100000000111010",
		342 => "1011111110001100",
		343 => "1011111011011111",
		344 => "1011111000110010",
		345 => "1011110110000110",
		346 => "1011110011011010",
		347 => "1011110000101111",
		348 => "1011101110000101",
		349 => "1011101011011100",
		350 => "1011101000110011",
		351 => "1011100110001011",
		352 => "1011100011100011",
		353 => "1011100000111100",
		354 => "1011011110010110",
		355 => "1011011011110001",
		356 => "1011011001001100",
		357 => "1011010110101000",
		358 => "1011010100000101",
		359 => "1011010001100010",
		360 => "1011001111000000",
		361 => "1011001100011111",
		362 => "1011001001111111",
		363 => "1011000111011111",
		364 => "1011000101000000",
		365 => "1011000010100010",
		366 => "1011000000000101",
		367 => "1010111101101000",
		368 => "1010111011001100",
		369 => "1010111000110001",
		370 => "1010110110010111",
		371 => "1010110011111110",
		372 => "1010110001100101",
		373 => "1010101111001101",
		374 => "1010101100110110",
		375 => "1010101010100000",
		376 => "1010101000001011",
		377 => "1010100101110110",
		378 => "1010100011100010",
		379 => "1010100001001111",
		380 => "1010011110111101",
		381 => "1010011100101100",
		382 => "1010011010011100",
		383 => "1010011000001100",
		384 => "1010010101111110",
		385 => "1010010011110000",
		386 => "1010010001100011",
		387 => "1010001111010111",
		388 => "1010001101001100",
		389 => "1010001011000010",
		390 => "1010001000111001",
		391 => "1010000110110000",
		392 => "1010000100101001",
		393 => "1010000010100010",
		394 => "1010000000011101",
		395 => "1001111110011000",
		396 => "1001111100010100",
		397 => "1001111010010001",
		398 => "1001111000001111",
		399 => "1001110110001110",
		400 => "1001110100001110",
		401 => "1001110010001111",
		402 => "1001110000010001",
		403 => "1001101110010100",
		404 => "1001101100011000",
		405 => "1001101010011101",
		406 => "1001101000100010",
		407 => "1001100110101001",
		408 => "1001100100110001",
		409 => "1001100010111010",
		410 => "1001100001000011",
		411 => "1001011111001110",
		412 => "1001011101011010",
		413 => "1001011011100110",
		414 => "1001011001110100",
		415 => "1001011000000011",
		416 => "1001010110010011",
		417 => "1001010100100100",
		418 => "1001010010110101",
		419 => "1001010001001000",
		420 => "1001001111011100",
		421 => "1001001101110001",
		422 => "1001001100000111",
		423 => "1001001010011110",
		424 => "1001001000110110",
		425 => "1001000111001111",
		426 => "1001000101101010",
		427 => "1001000100000101",
		428 => "1001000010100001",
		429 => "1001000000111111",
		430 => "1000111111011101",
		431 => "1000111101111101",
		432 => "1000111100011110",
		433 => "1000111010111111",
		434 => "1000111001100010",
		435 => "1000111000000110",
		436 => "1000110110101011",
		437 => "1000110101010001",
		438 => "1000110011111001",
		439 => "1000110010100001",
		440 => "1000110001001010",
		441 => "1000101111110101",
		442 => "1000101110100001",
		443 => "1000101101001110",
		444 => "1000101011111100",
		445 => "1000101010101011",
		446 => "1000101001011011",
		447 => "1000101000001100",
		448 => "1000100110111111",
		449 => "1000100101110010",
		450 => "1000100100100111",
		451 => "1000100011011101",
		452 => "1000100010010100",
		453 => "1000100001001100",
		454 => "1000100000000110",
		455 => "1000011111000000",
		456 => "1000011101111100",
		457 => "1000011100111001",
		458 => "1000011011110111",
		459 => "1000011010110110",
		460 => "1000011001110110",
		461 => "1000011000111000",
		462 => "1000010111111011",
		463 => "1000010110111110",
		464 => "1000010110000011",
		465 => "1000010101001010",
		466 => "1000010100010001",
		467 => "1000010011011010",
		468 => "1000010010100011",
		469 => "1000010001101110",
		470 => "1000010000111011",
		471 => "1000010000001000",
		472 => "1000001111010110",
		473 => "1000001110100110",
		474 => "1000001101110111",
		475 => "1000001101001001",
		476 => "1000001100011101",
		477 => "1000001011110001",
		478 => "1000001011000111",
		479 => "1000001010011110",
		480 => "1000001001110110",
		481 => "1000001001001111",
		482 => "1000001000101010",
		483 => "1000001000000110",
		484 => "1000000111100011",
		485 => "1000000111000001",
		486 => "1000000110100001",
		487 => "1000000110000001",
		488 => "1000000101100011",
		489 => "1000000101000110",
		490 => "1000000100101011",
		491 => "1000000100010000",
		492 => "1000000011110111",
		493 => "1000000011011111",
		494 => "1000000011001000",
		495 => "1000000010110011",
		496 => "1000000010011110",
		497 => "1000000010001011",
		498 => "1000000001111001",
		499 => "1000000001101001",
		500 => "1000000001011001",
		501 => "1000000001001011",
		502 => "1000000000111110",
		503 => "1000000000110010",
		504 => "1000000000101000",
		505 => "1000000000011111",
		506 => "1000000000010111",
		507 => "1000000000010000",
		508 => "1000000000001010",
		509 => "1000000000000110",
		510 => "1000000000000011",
		511 => "1000000000000001"
		);

	constant im_64: arr := (
		0 => "0000000000000000",
		1 => "0000000011001001",
		2 => "0000000110010010",
		3 => "0000001001011011",
		4 => "0000001100100100",
		5 => "0000001111101101",
		6 => "0000010010110110",
		7 => "0000010101111110",
		8 => "0000011001000111",
		9 => "0000011100010000",
		10 => "0000011111011001",
		11 => "0000100010100001",
		12 => "0000100101101010",
		13 => "0000101000110010",
		14 => "0000101011111011",
		15 => "0000101111000011",
		16 => "0000110010001011",
		17 => "0000110101010011",
		18 => "0000111000011011",
		19 => "0000111011100011",
		20 => "0000111110101011",
		21 => "0001000001110010",
		22 => "0001000100111001",
		23 => "0001001000000000",
		24 => "0001001011000111",
		25 => "0001001110001110",
		26 => "0001010001010101",
		27 => "0001010100011011",
		28 => "0001010111100001",
		29 => "0001011010100111",
		30 => "0001011101101101",
		31 => "0001100000110011",
		32 => "0001100011111000",
		33 => "0001100110111101",
		34 => "0001101010000010",
		35 => "0001101101000110",
		36 => "0001110000001011",
		37 => "0001110011001111",
		38 => "0001110110010011",
		39 => "0001111001010110",
		40 => "0001111100011001",
		41 => "0001111111011100",
		42 => "0010000010011111",
		43 => "0010000101100001",
		44 => "0010001000100011",
		45 => "0010001011100100",
		46 => "0010001110100110",
		47 => "0010010001100111",
		48 => "0010010100100111",
		49 => "0010010111100111",
		50 => "0010011010100111",
		51 => "0010011101100111",
		52 => "0010100000100110",
		53 => "0010100011100101",
		54 => "0010100110100011",
		55 => "0010101001100001",
		56 => "0010101100011110",
		57 => "0010101111011011",
		58 => "0010110010011000",
		59 => "0010110101010100",
		60 => "0010111000010000",
		61 => "0010111011001100",
		62 => "0010111110000110",
		63 => "0011000001000001",
		64 => "0011000011111011",
		65 => "0011000110110100",
		66 => "0011001001101101",
		67 => "0011001100100110",
		68 => "0011001111011110",
		69 => "0011010010010110",
		70 => "0011010101001101",
		71 => "0011011000000011",
		72 => "0011011010111001",
		73 => "0011011101101111",
		74 => "0011100000100100",
		75 => "0011100011011000",
		76 => "0011100110001100",
		77 => "0011101000111111",
		78 => "0011101011110010",
		79 => "0011101110100100",
		80 => "0011110001010110",
		81 => "0011110100000111",
		82 => "0011110110110111",
		83 => "0011111001100111",
		84 => "0011111100010110",
		85 => "0011111111000101",
		86 => "0100000001110011",
		87 => "0100000100100000",
		88 => "0100000111001101",
		89 => "0100001001111001",
		90 => "0100001100100101",
		91 => "0100001111010000",
		92 => "0100010001111010",
		93 => "0100010100100011",
		94 => "0100010111001100",
		95 => "0100011001110100",
		96 => "0100011100011100",
		97 => "0100011111000011",
		98 => "0100100001101001",
		99 => "0100100100001110",
		100 => "0100100110110011",
		101 => "0100101001010111",
		102 => "0100101011111010",
		103 => "0100101110011101",
		104 => "0100110000111111",
		105 => "0100110011100000",
		106 => "0100110110000000",
		107 => "0100111000100000",
		108 => "0100111010111111",
		109 => "0100111101011101",
		110 => "0100111111111010",
		111 => "0101000010010111",
		112 => "0101000100110011",
		113 => "0101000111001110",
		114 => "0101001001101000",
		115 => "0101001100000001",
		116 => "0101001110011010",
		117 => "0101010000110010",
		118 => "0101010011001001",
		119 => "0101010101011111",
		120 => "0101010111110100",
		121 => "0101011010001001",
		122 => "0101011100011101",
		123 => "0101011110110000",
		124 => "0101100001000010",
		125 => "0101100011010011",
		126 => "0101100101100011",
		127 => "0101100111110011",
		128 => "0101101010000001",
		129 => "0101101100001111",
		130 => "0101101110011100",
		131 => "0101110000101000",
		132 => "0101110010110011",
		133 => "0101110100111101",
		134 => "0101110111000110",
		135 => "0101111001001111",
		136 => "0101111011010110",
		137 => "0101111101011101",
		138 => "0101111111100010",
		139 => "0110000001100111",
		140 => "0110000011101011",
		141 => "0110000101101110",
		142 => "0110000111110000",
		143 => "0110001001110001",
		144 => "0110001011110001",
		145 => "0110001101110000",
		146 => "0110001111101110",
		147 => "0110010001101011",
		148 => "0110010011100111",
		149 => "0110010101100010",
		150 => "0110010111011101",
		151 => "0110011001010110",
		152 => "0110011011001110",
		153 => "0110011101000101",
		154 => "0110011110111100",
		155 => "0110100000110001",
		156 => "0110100010100101",
		157 => "0110100100011001",
		158 => "0110100110001011",
		159 => "0110100111111100",
		160 => "0110101001101100",
		161 => "0110101011011011",
		162 => "0110101101001010",
		163 => "0110101110110111",
		164 => "0110110000100011",
		165 => "0110110010001110",
		166 => "0110110011111000",
		167 => "0110110101100001",
		168 => "0110110111001001",
		169 => "0110111000110000",
		170 => "0110111010010101",
		171 => "0110111011111010",
		172 => "0110111101011110",
		173 => "0110111111000000",
		174 => "0111000000100010",
		175 => "0111000010000010",
		176 => "0111000011100001",
		177 => "0111000101000000",
		178 => "0111000110011101",
		179 => "0111000111111001",
		180 => "0111001001010100",
		181 => "0111001010101110",
		182 => "0111001100000110",
		183 => "0111001101011110",
		184 => "0111001110110101",
		185 => "0111010000001010",
		186 => "0111010001011110",
		187 => "0111010010110001",
		188 => "0111010100000011",
		189 => "0111010101010100",
		190 => "0111010110100100",
		191 => "0111010111110011",
		192 => "0111011001000000",
		193 => "0111011010001101",
		194 => "0111011011011000",
		195 => "0111011100100010",
		196 => "0111011101101011",
		197 => "0111011110110011",
		198 => "0111011111111001",
		199 => "0111100000111111",
		200 => "0111100010000011",
		201 => "0111100011000110",
		202 => "0111100100001000",
		203 => "0111100101001001",
		204 => "0111100110001001",
		205 => "0111100111000111",
		206 => "0111101000000100",
		207 => "0111101001000001",
		208 => "0111101001111100",
		209 => "0111101010110101",
		210 => "0111101011101110",
		211 => "0111101100100101",
		212 => "0111101101011100",
		213 => "0111101110010001",
		214 => "0111101111000100",
		215 => "0111101111110111",
		216 => "0111110000101001",
		217 => "0111110001011001",
		218 => "0111110010001000",
		219 => "0111110010110110",
		220 => "0111110011100010",
		221 => "0111110100001110",
		222 => "0111110100111000",
		223 => "0111110101100001",
		224 => "0111110110001001",
		225 => "0111110110110000",
		226 => "0111110111010101",
		227 => "0111110111111001",
		228 => "0111111000011100",
		229 => "0111111000111110",
		230 => "0111111001011110",
		231 => "0111111001111110",
		232 => "0111111010011100",
		233 => "0111111010111001",
		234 => "0111111011010100",
		235 => "0111111011101111",
		236 => "0111111100001000",
		237 => "0111111100100000",
		238 => "0111111100110111",
		239 => "0111111101001100",
		240 => "0111111101100001",
		241 => "0111111101110100",
		242 => "0111111110000110",
		243 => "0111111110010110",
		244 => "0111111110100110",
		245 => "0111111110110100",
		246 => "0111111111000001",
		247 => "0111111111001101",
		248 => "0111111111010111",
		249 => "0111111111100000",
		250 => "0111111111101000",
		251 => "0111111111101111",
		252 => "0111111111110101",
		253 => "0111111111111001",
		254 => "0111111111111100",
		255 => "0111111111111110",
		256 => "0111111111111111",
		257 => "0111111111111110",
		258 => "0111111111111100",
		259 => "0111111111111001",
		260 => "0111111111110101",
		261 => "0111111111101111",
		262 => "0111111111101000",
		263 => "0111111111100000",
		264 => "0111111111010111",
		265 => "0111111111001101",
		266 => "0111111111000001",
		267 => "0111111110110100",
		268 => "0111111110100110",
		269 => "0111111110010110",
		270 => "0111111110000110",
		271 => "0111111101110100",
		272 => "0111111101100001",
		273 => "0111111101001100",
		274 => "0111111100110111",
		275 => "0111111100100000",
		276 => "0111111100001000",
		277 => "0111111011101111",
		278 => "0111111011010100",
		279 => "0111111010111001",
		280 => "0111111010011100",
		281 => "0111111001111110",
		282 => "0111111001011110",
		283 => "0111111000111110",
		284 => "0111111000011100",
		285 => "0111110111111001",
		286 => "0111110111010101",
		287 => "0111110110110000",
		288 => "0111110110001001",
		289 => "0111110101100001",
		290 => "0111110100111000",
		291 => "0111110100001110",
		292 => "0111110011100010",
		293 => "0111110010110110",
		294 => "0111110010001000",
		295 => "0111110001011001",
		296 => "0111110000101001",
		297 => "0111101111110111",
		298 => "0111101111000100",
		299 => "0111101110010001",
		300 => "0111101101011100",
		301 => "0111101100100101",
		302 => "0111101011101110",
		303 => "0111101010110101",
		304 => "0111101001111100",
		305 => "0111101001000001",
		306 => "0111101000000100",
		307 => "0111100111000111",
		308 => "0111100110001001",
		309 => "0111100101001001",
		310 => "0111100100001000",
		311 => "0111100011000110",
		312 => "0111100010000011",
		313 => "0111100000111111",
		314 => "0111011111111001",
		315 => "0111011110110011",
		316 => "0111011101101011",
		317 => "0111011100100010",
		318 => "0111011011011000",
		319 => "0111011010001101",
		320 => "0111011001000000",
		321 => "0111010111110011",
		322 => "0111010110100100",
		323 => "0111010101010100",
		324 => "0111010100000011",
		325 => "0111010010110001",
		326 => "0111010001011110",
		327 => "0111010000001010",
		328 => "0111001110110101",
		329 => "0111001101011110",
		330 => "0111001100000110",
		331 => "0111001010101110",
		332 => "0111001001010100",
		333 => "0111000111111001",
		334 => "0111000110011101",
		335 => "0111000101000000",
		336 => "0111000011100001",
		337 => "0111000010000010",
		338 => "0111000000100010",
		339 => "0110111111000000",
		340 => "0110111101011110",
		341 => "0110111011111010",
		342 => "0110111010010101",
		343 => "0110111000110000",
		344 => "0110110111001001",
		345 => "0110110101100001",
		346 => "0110110011111000",
		347 => "0110110010001110",
		348 => "0110110000100011",
		349 => "0110101110110111",
		350 => "0110101101001010",
		351 => "0110101011011011",
		352 => "0110101001101100",
		353 => "0110100111111100",
		354 => "0110100110001011",
		355 => "0110100100011001",
		356 => "0110100010100101",
		357 => "0110100000110001",
		358 => "0110011110111100",
		359 => "0110011101000101",
		360 => "0110011011001110",
		361 => "0110011001010110",
		362 => "0110010111011101",
		363 => "0110010101100010",
		364 => "0110010011100111",
		365 => "0110010001101011",
		366 => "0110001111101110",
		367 => "0110001101110000",
		368 => "0110001011110001",
		369 => "0110001001110001",
		370 => "0110000111110000",
		371 => "0110000101101110",
		372 => "0110000011101011",
		373 => "0110000001100111",
		374 => "0101111111100010",
		375 => "0101111101011101",
		376 => "0101111011010110",
		377 => "0101111001001111",
		378 => "0101110111000110",
		379 => "0101110100111101",
		380 => "0101110010110011",
		381 => "0101110000101000",
		382 => "0101101110011100",
		383 => "0101101100001111",
		384 => "0101101010000001",
		385 => "0101100111110011",
		386 => "0101100101100011",
		387 => "0101100011010011",
		388 => "0101100001000010",
		389 => "0101011110110000",
		390 => "0101011100011101",
		391 => "0101011010001001",
		392 => "0101010111110100",
		393 => "0101010101011111",
		394 => "0101010011001001",
		395 => "0101010000110010",
		396 => "0101001110011010",
		397 => "0101001100000001",
		398 => "0101001001101000",
		399 => "0101000111001110",
		400 => "0101000100110011",
		401 => "0101000010010111",
		402 => "0100111111111010",
		403 => "0100111101011101",
		404 => "0100111010111111",
		405 => "0100111000100000",
		406 => "0100110110000000",
		407 => "0100110011100000",
		408 => "0100110000111111",
		409 => "0100101110011101",
		410 => "0100101011111010",
		411 => "0100101001010111",
		412 => "0100100110110011",
		413 => "0100100100001110",
		414 => "0100100001101001",
		415 => "0100011111000011",
		416 => "0100011100011100",
		417 => "0100011001110100",
		418 => "0100010111001100",
		419 => "0100010100100011",
		420 => "0100010001111010",
		421 => "0100001111010000",
		422 => "0100001100100101",
		423 => "0100001001111001",
		424 => "0100000111001101",
		425 => "0100000100100000",
		426 => "0100000001110011",
		427 => "0011111111000101",
		428 => "0011111100010110",
		429 => "0011111001100111",
		430 => "0011110110110111",
		431 => "0011110100000111",
		432 => "0011110001010110",
		433 => "0011101110100100",
		434 => "0011101011110010",
		435 => "0011101000111111",
		436 => "0011100110001100",
		437 => "0011100011011000",
		438 => "0011100000100100",
		439 => "0011011101101111",
		440 => "0011011010111001",
		441 => "0011011000000011",
		442 => "0011010101001101",
		443 => "0011010010010110",
		444 => "0011001111011110",
		445 => "0011001100100110",
		446 => "0011001001101101",
		447 => "0011000110110100",
		448 => "0011000011111011",
		449 => "0011000001000001",
		450 => "0010111110000110",
		451 => "0010111011001100",
		452 => "0010111000010000",
		453 => "0010110101010100",
		454 => "0010110010011000",
		455 => "0010101111011011",
		456 => "0010101100011110",
		457 => "0010101001100001",
		458 => "0010100110100011",
		459 => "0010100011100101",
		460 => "0010100000100110",
		461 => "0010011101100111",
		462 => "0010011010100111",
		463 => "0010010111100111",
		464 => "0010010100100111",
		465 => "0010010001100111",
		466 => "0010001110100110",
		467 => "0010001011100100",
		468 => "0010001000100011",
		469 => "0010000101100001",
		470 => "0010000010011111",
		471 => "0001111111011100",
		472 => "0001111100011001",
		473 => "0001111001010110",
		474 => "0001110110010011",
		475 => "0001110011001111",
		476 => "0001110000001011",
		477 => "0001101101000110",
		478 => "0001101010000010",
		479 => "0001100110111101",
		480 => "0001100011111000",
		481 => "0001100000110011",
		482 => "0001011101101101",
		483 => "0001011010100111",
		484 => "0001010111100001",
		485 => "0001010100011011",
		486 => "0001010001010101",
		487 => "0001001110001110",
		488 => "0001001011000111",
		489 => "0001001000000000",
		490 => "0001000100111001",
		491 => "0001000001110010",
		492 => "0000111110101011",
		493 => "0000111011100011",
		494 => "0000111000011011",
		495 => "0000110101010011",
		496 => "0000110010001011",
		497 => "0000101111000011",
		498 => "0000101011111011",
		499 => "0000101000110010",
		500 => "0000100101101010",
		501 => "0000100010100001",
		502 => "0000011111011001",
		503 => "0000011100010000",
		504 => "0000011001000111",
		505 => "0000010101111110",
		506 => "0000010010110110",
		507 => "0000001111101101",
		508 => "0000001100100100",
		509 => "0000001001011011",
		510 => "0000000110010010",
		511 => "0000000011001001"
		);
end;
