library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fft_twiddle_factors_64 is
	constant tw_size:           integer := 14;
	constant tw_array_size_exp: integer := 6;
	
	type arr is array (0 to 2**(tw_array_size_exp - 1) - 1) of signed(tw_size - 1 downto 0);

	constant re_64: arr := (
		0 => "01111111111111",
		1 => "01111111010111",
		2 => "01111101100001",
		3 => "01111010011110",
		4 => "01110110001111",
		5 => "01110000110111",
		6 => "01101010011010",
		7 => "01100010111011",
		8 => "01011010011111",
		9 => "01010001001100",
		10 => "01000111000110",
		11 => "00111100010101",
		12 => "00110000111110",
		13 => "00100101001001",
		14 => "00011000111101",
		15 => "00001100100010",
		16 => "00000000000000",
		17 => "11110011011101",
		18 => "11100111000010",
		19 => "11011010110110",
		20 => "11001111000001",
		21 => "11000011101010",
		22 => "10111000111001",
		23 => "10101110110011",
		24 => "10100101100000",
		25 => "10011101000100",
		26 => "10010101100101",
		27 => "10001111001000",
		28 => "10001001110000",
		29 => "10000101100001",
		30 => "10000010011110",
		31 => "10000000101000"
		);

	constant im_64: arr := (
		0 => "00000000000000",
		1 => "00001100100010",
		2 => "00011000111101",
		3 => "00100101001001",
		4 => "00110000111110",
		5 => "00111100010101",
		6 => "01000111000110",
		7 => "01010001001100",
		8 => "01011010011111",
		9 => "01100010111011",
		10 => "01101010011010",
		11 => "01110000110111",
		12 => "01110110001111",
		13 => "01111010011110",
		14 => "01111101100001",
		15 => "01111111010111",
		16 => "01111111111111",
		17 => "01111111010111",
		18 => "01111101100001",
		19 => "01111010011110",
		20 => "01110110001111",
		21 => "01110000110111",
		22 => "01101010011010",
		23 => "01100010111011",
		24 => "01011010011111",
		25 => "01010001001100",
		26 => "01000111000110",
		27 => "00111100010101",
		28 => "00110000111110",
		29 => "00100101001001",
		30 => "00011000111101",
		31 => "00001100100010"
		);
end;
