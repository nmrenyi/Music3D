library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package trans_pkg is
    type cube_vector is array(7 downto 0) of std_logic_vector(63 downto 0);
end package;